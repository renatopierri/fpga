module shifter(
	input [7:0] inp,			
	input [1:0] shift_cntrl,	
	output reg [15:0] shift_out
);
 
	// Tornando todas entradas sensíveis ao evento:
	always@(inp, shift_cntrl) begin
		if (shift_cntrl == 2'b01)
			shift_out = (inp << 4);
		else if (shift_cntrl == 2'b10)
			shift_out = (inp << 8);
		else
			shift_out = inp;
	end
endmodule 